module SmallCircle(output Ci, input Gi);
  
 // buf  (Ci, Gi);
    assign Ci=Gi;
  
endmodule
